// hps.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module hps (
		input  wire [15:0] arduino_io_external_connection_in_port,  // arduino_io_external_connection.in_port
		output wire [15:0] arduino_io_external_connection_out_port, //                               .out_port
		input  wire        clk_clk,                                 //                            clk.clk
		input  wire [31:0] gpio0_external_connection_in_port,       //      gpio0_external_connection.in_port
		output wire [31:0] gpio0_external_connection_out_port,      //                               .out_port
		input  wire [31:0] gpio1_external_connection_in_port,       //      gpio1_external_connection.in_port
		output wire [31:0] gpio1_external_connection_out_port,      //                               .out_port
		inout  wire        hps_io_hps_io_sdio_inst_CMD,             //                         hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,              //                               .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,              //                               .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,             //                               .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,              //                               .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,              //                               .hps_io_sdio_inst_D3
		input  wire        hps_io_hps_io_uart0_inst_RX,             //                               .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,             //                               .hps_io_uart0_inst_TX
		input  wire [1:0]  keys_external_connection_export,         //       keys_external_connection.export
		output wire [7:0]  led_external_connection_export,          //        led_external_connection.export
		output wire [12:0] memory_mem_a,                            //                         memory.mem_a
		output wire [2:0]  memory_mem_ba,                           //                               .mem_ba
		output wire        memory_mem_ck,                           //                               .mem_ck
		output wire        memory_mem_ck_n,                         //                               .mem_ck_n
		output wire        memory_mem_cke,                          //                               .mem_cke
		output wire        memory_mem_cs_n,                         //                               .mem_cs_n
		output wire        memory_mem_ras_n,                        //                               .mem_ras_n
		output wire        memory_mem_cas_n,                        //                               .mem_cas_n
		output wire        memory_mem_we_n,                         //                               .mem_we_n
		output wire        memory_mem_reset_n,                      //                               .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                           //                               .mem_dq
		inout  wire        memory_mem_dqs,                          //                               .mem_dqs
		inout  wire			 memory_mem_dqs_n,                        //                               .mem_dqs_n
		output wire        memory_mem_odt,                          //                               .mem_odt
		output wire        memory_mem_dm,                           //                               .mem_dm
		input  wire        memory_oct_rzqin,                        //                               .oct_rzqin
		input  wire [3:0]  sw_external_connection_export            //         sw_external_connection.export
	);

	wire         hps_h2f_reset_reset;                        // HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire   [1:0] hps_h2f_lw_axi_master_awburst;              // HPS:h2f_lw_AWBURST -> mm_interconnect_0:HPS_h2f_lw_axi_master_awburst
	wire   [3:0] hps_h2f_lw_axi_master_arlen;                // HPS:h2f_lw_ARLEN -> mm_interconnect_0:HPS_h2f_lw_axi_master_arlen
	wire   [3:0] hps_h2f_lw_axi_master_wstrb;                // HPS:h2f_lw_WSTRB -> mm_interconnect_0:HPS_h2f_lw_axi_master_wstrb
	wire         hps_h2f_lw_axi_master_wready;               // mm_interconnect_0:HPS_h2f_lw_axi_master_wready -> HPS:h2f_lw_WREADY
	wire  [11:0] hps_h2f_lw_axi_master_rid;                  // mm_interconnect_0:HPS_h2f_lw_axi_master_rid -> HPS:h2f_lw_RID
	wire         hps_h2f_lw_axi_master_rready;               // HPS:h2f_lw_RREADY -> mm_interconnect_0:HPS_h2f_lw_axi_master_rready
	wire   [3:0] hps_h2f_lw_axi_master_awlen;                // HPS:h2f_lw_AWLEN -> mm_interconnect_0:HPS_h2f_lw_axi_master_awlen
	wire  [11:0] hps_h2f_lw_axi_master_wid;                  // HPS:h2f_lw_WID -> mm_interconnect_0:HPS_h2f_lw_axi_master_wid
	wire   [3:0] hps_h2f_lw_axi_master_arcache;              // HPS:h2f_lw_ARCACHE -> mm_interconnect_0:HPS_h2f_lw_axi_master_arcache
	wire         hps_h2f_lw_axi_master_wvalid;               // HPS:h2f_lw_WVALID -> mm_interconnect_0:HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_h2f_lw_axi_master_araddr;               // HPS:h2f_lw_ARADDR -> mm_interconnect_0:HPS_h2f_lw_axi_master_araddr
	wire   [2:0] hps_h2f_lw_axi_master_arprot;               // HPS:h2f_lw_ARPROT -> mm_interconnect_0:HPS_h2f_lw_axi_master_arprot
	wire   [2:0] hps_h2f_lw_axi_master_awprot;               // HPS:h2f_lw_AWPROT -> mm_interconnect_0:HPS_h2f_lw_axi_master_awprot
	wire  [31:0] hps_h2f_lw_axi_master_wdata;                // HPS:h2f_lw_WDATA -> mm_interconnect_0:HPS_h2f_lw_axi_master_wdata
	wire         hps_h2f_lw_axi_master_arvalid;              // HPS:h2f_lw_ARVALID -> mm_interconnect_0:HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_h2f_lw_axi_master_awcache;              // HPS:h2f_lw_AWCACHE -> mm_interconnect_0:HPS_h2f_lw_axi_master_awcache
	wire  [11:0] hps_h2f_lw_axi_master_arid;                 // HPS:h2f_lw_ARID -> mm_interconnect_0:HPS_h2f_lw_axi_master_arid
	wire   [1:0] hps_h2f_lw_axi_master_arlock;               // HPS:h2f_lw_ARLOCK -> mm_interconnect_0:HPS_h2f_lw_axi_master_arlock
	wire   [1:0] hps_h2f_lw_axi_master_awlock;               // HPS:h2f_lw_AWLOCK -> mm_interconnect_0:HPS_h2f_lw_axi_master_awlock
	wire  [20:0] hps_h2f_lw_axi_master_awaddr;               // HPS:h2f_lw_AWADDR -> mm_interconnect_0:HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_h2f_lw_axi_master_bresp;                // mm_interconnect_0:HPS_h2f_lw_axi_master_bresp -> HPS:h2f_lw_BRESP
	wire         hps_h2f_lw_axi_master_arready;              // mm_interconnect_0:HPS_h2f_lw_axi_master_arready -> HPS:h2f_lw_ARREADY
	wire  [31:0] hps_h2f_lw_axi_master_rdata;                // mm_interconnect_0:HPS_h2f_lw_axi_master_rdata -> HPS:h2f_lw_RDATA
	wire         hps_h2f_lw_axi_master_awready;              // mm_interconnect_0:HPS_h2f_lw_axi_master_awready -> HPS:h2f_lw_AWREADY
	wire   [1:0] hps_h2f_lw_axi_master_arburst;              // HPS:h2f_lw_ARBURST -> mm_interconnect_0:HPS_h2f_lw_axi_master_arburst
	wire   [2:0] hps_h2f_lw_axi_master_arsize;               // HPS:h2f_lw_ARSIZE -> mm_interconnect_0:HPS_h2f_lw_axi_master_arsize
	wire         hps_h2f_lw_axi_master_bready;               // HPS:h2f_lw_BREADY -> mm_interconnect_0:HPS_h2f_lw_axi_master_bready
	wire         hps_h2f_lw_axi_master_rlast;                // mm_interconnect_0:HPS_h2f_lw_axi_master_rlast -> HPS:h2f_lw_RLAST
	wire         hps_h2f_lw_axi_master_wlast;                // HPS:h2f_lw_WLAST -> mm_interconnect_0:HPS_h2f_lw_axi_master_wlast
	wire   [1:0] hps_h2f_lw_axi_master_rresp;                // mm_interconnect_0:HPS_h2f_lw_axi_master_rresp -> HPS:h2f_lw_RRESP
	wire  [11:0] hps_h2f_lw_axi_master_awid;                 // HPS:h2f_lw_AWID -> mm_interconnect_0:HPS_h2f_lw_axi_master_awid
	wire  [11:0] hps_h2f_lw_axi_master_bid;                  // mm_interconnect_0:HPS_h2f_lw_axi_master_bid -> HPS:h2f_lw_BID
	wire         hps_h2f_lw_axi_master_bvalid;               // mm_interconnect_0:HPS_h2f_lw_axi_master_bvalid -> HPS:h2f_lw_BVALID
	wire   [2:0] hps_h2f_lw_axi_master_awsize;               // HPS:h2f_lw_AWSIZE -> mm_interconnect_0:HPS_h2f_lw_axi_master_awsize
	wire         hps_h2f_lw_axi_master_awvalid;              // HPS:h2f_lw_AWVALID -> mm_interconnect_0:HPS_h2f_lw_axi_master_awvalid
	wire         hps_h2f_lw_axi_master_rvalid;               // mm_interconnect_0:HPS_h2f_lw_axi_master_rvalid -> HPS:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;         // keys:readdata -> mm_interconnect_0:keys_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;          // mm_interconnect_0:keys_s1_address -> keys:address
	wire         mm_interconnect_0_led_s1_chipselect;        // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;          // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;           // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;             // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;         // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;           // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;            // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_gpio0_s1_chipselect;      // mm_interconnect_0:gpio0_s1_chipselect -> gpio0:chipselect
	wire  [31:0] mm_interconnect_0_gpio0_s1_readdata;        // gpio0:readdata -> mm_interconnect_0:gpio0_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio0_s1_address;         // mm_interconnect_0:gpio0_s1_address -> gpio0:address
	wire         mm_interconnect_0_gpio0_s1_write;           // mm_interconnect_0:gpio0_s1_write -> gpio0:write_n
	wire  [31:0] mm_interconnect_0_gpio0_s1_writedata;       // mm_interconnect_0:gpio0_s1_writedata -> gpio0:writedata
	wire         mm_interconnect_0_gpio1_s1_chipselect;      // mm_interconnect_0:gpio1_s1_chipselect -> gpio1:chipselect
	wire  [31:0] mm_interconnect_0_gpio1_s1_readdata;        // gpio1:readdata -> mm_interconnect_0:gpio1_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio1_s1_address;         // mm_interconnect_0:gpio1_s1_address -> gpio1:address
	wire         mm_interconnect_0_gpio1_s1_write;           // mm_interconnect_0:gpio1_s1_write -> gpio1:write_n
	wire  [31:0] mm_interconnect_0_gpio1_s1_writedata;       // mm_interconnect_0:gpio1_s1_writedata -> gpio1:writedata
	wire         mm_interconnect_0_arduino_io_s1_chipselect; // mm_interconnect_0:Arduino_io_s1_chipselect -> Arduino_io:chipselect
	wire  [31:0] mm_interconnect_0_arduino_io_s1_readdata;   // Arduino_io:readdata -> mm_interconnect_0:Arduino_io_s1_readdata
	wire   [1:0] mm_interconnect_0_arduino_io_s1_address;    // mm_interconnect_0:Arduino_io_s1_address -> Arduino_io:address
	wire         mm_interconnect_0_arduino_io_s1_write;      // mm_interconnect_0:Arduino_io_s1_write -> Arduino_io:write_n
	wire  [31:0] mm_interconnect_0_arduino_io_s1_writedata;  // mm_interconnect_0:Arduino_io_s1_writedata -> Arduino_io:writedata
	wire         rst_controller_reset_out_reset;             // rst_controller:reset_out -> [Arduino_io:reset_n, gpio0:reset_n, gpio1:reset_n, keys:reset_n, led:reset_n, mm_interconnect_0:keys_reset_reset_bridge_in_reset_reset, sw:reset_n]
	wire         rst_controller_001_reset_out_reset;         // rst_controller_001:reset_out -> mm_interconnect_0:HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	hps_Arduino_io arduino_io (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_arduino_io_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_arduino_io_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_arduino_io_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_arduino_io_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_arduino_io_s1_readdata),   //                    .readdata
		.in_port    (arduino_io_external_connection_in_port),     // external_connection.export
		.out_port   (arduino_io_external_connection_out_port)     //                    .export
	);

	hps_HPS #(
		.F2S_Width (1),
		.S2F_Width (1)
	) hps (
		.mem_a                (memory_mem_a),                  //            memory.mem_a
		.mem_ba               (memory_mem_ba),                 //                  .mem_ba
		.mem_ck               (memory_mem_ck),                 //                  .mem_ck
		.mem_ck_n             (memory_mem_ck_n),               //                  .mem_ck_n
		.mem_cke              (memory_mem_cke),                //                  .mem_cke
		.mem_cs_n             (memory_mem_cs_n),               //                  .mem_cs_n
		.mem_ras_n            (memory_mem_ras_n),              //                  .mem_ras_n
		.mem_cas_n            (memory_mem_cas_n),              //                  .mem_cas_n
		.mem_we_n             (memory_mem_we_n),               //                  .mem_we_n
		.mem_reset_n          (memory_mem_reset_n),            //                  .mem_reset_n
		.mem_dq               (memory_mem_dq),                 //                  .mem_dq
		.mem_dqs              (memory_mem_dqs),                //                  .mem_dqs
		.mem_dqs_n            (memory_mem_dqs_n),              //                  .mem_dqs_n
		.mem_odt              (memory_mem_odt),                //                  .mem_odt
		.mem_dm               (memory_mem_dm),                 //                  .mem_dm
		.oct_rzqin            (memory_oct_rzqin),              //                  .oct_rzqin
		.hps_io_sdio_inst_CMD (hps_io_hps_io_sdio_inst_CMD),   //            hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0  (hps_io_hps_io_sdio_inst_D0),    //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1  (hps_io_hps_io_sdio_inst_D1),    //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK (hps_io_hps_io_sdio_inst_CLK),   //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2  (hps_io_hps_io_sdio_inst_D2),    //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3  (hps_io_hps_io_sdio_inst_D3),    //                  .hps_io_sdio_inst_D3
		.hps_io_uart0_inst_RX (hps_io_hps_io_uart0_inst_RX),   //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX (hps_io_hps_io_uart0_inst_TX),   //                  .hps_io_uart0_inst_TX
		.h2f_rst_n            (hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk          (clk_clk),                       //     h2f_axi_clock.clk
		.h2f_AWID             (),                              //    h2f_axi_master.awid
		.h2f_AWADDR           (),                              //                  .awaddr
		.h2f_AWLEN            (),                              //                  .awlen
		.h2f_AWSIZE           (),                              //                  .awsize
		.h2f_AWBURST          (),                              //                  .awburst
		.h2f_AWLOCK           (),                              //                  .awlock
		.h2f_AWCACHE          (),                              //                  .awcache
		.h2f_AWPROT           (),                              //                  .awprot
		.h2f_AWVALID          (),                              //                  .awvalid
		.h2f_AWREADY          (),                              //                  .awready
		.h2f_WID              (),                              //                  .wid
		.h2f_WDATA            (),                              //                  .wdata
		.h2f_WSTRB            (),                              //                  .wstrb
		.h2f_WLAST            (),                              //                  .wlast
		.h2f_WVALID           (),                              //                  .wvalid
		.h2f_WREADY           (),                              //                  .wready
		.h2f_BID              (),                              //                  .bid
		.h2f_BRESP            (),                              //                  .bresp
		.h2f_BVALID           (),                              //                  .bvalid
		.h2f_BREADY           (),                              //                  .bready
		.h2f_ARID             (),                              //                  .arid
		.h2f_ARADDR           (),                              //                  .araddr
		.h2f_ARLEN            (),                              //                  .arlen
		.h2f_ARSIZE           (),                              //                  .arsize
		.h2f_ARBURST          (),                              //                  .arburst
		.h2f_ARLOCK           (),                              //                  .arlock
		.h2f_ARCACHE          (),                              //                  .arcache
		.h2f_ARPROT           (),                              //                  .arprot
		.h2f_ARVALID          (),                              //                  .arvalid
		.h2f_ARREADY          (),                              //                  .arready
		.h2f_RID              (),                              //                  .rid
		.h2f_RDATA            (),                              //                  .rdata
		.h2f_RRESP            (),                              //                  .rresp
		.h2f_RLAST            (),                              //                  .rlast
		.h2f_RVALID           (),                              //                  .rvalid
		.h2f_RREADY           (),                              //                  .rready
		.f2h_axi_clk          (clk_clk),                       //     f2h_axi_clock.clk
		.f2h_AWID             (),                              //     f2h_axi_slave.awid
		.f2h_AWADDR           (),                              //                  .awaddr
		.f2h_AWLEN            (),                              //                  .awlen
		.f2h_AWSIZE           (),                              //                  .awsize
		.f2h_AWBURST          (),                              //                  .awburst
		.f2h_AWLOCK           (),                              //                  .awlock
		.f2h_AWCACHE          (),                              //                  .awcache
		.f2h_AWPROT           (),                              //                  .awprot
		.f2h_AWVALID          (),                              //                  .awvalid
		.f2h_AWREADY          (),                              //                  .awready
		.f2h_AWUSER           (),                              //                  .awuser
		.f2h_WID              (),                              //                  .wid
		.f2h_WDATA            (),                              //                  .wdata
		.f2h_WSTRB            (),                              //                  .wstrb
		.f2h_WLAST            (),                              //                  .wlast
		.f2h_WVALID           (),                              //                  .wvalid
		.f2h_WREADY           (),                              //                  .wready
		.f2h_BID              (),                              //                  .bid
		.f2h_BRESP            (),                              //                  .bresp
		.f2h_BVALID           (),                              //                  .bvalid
		.f2h_BREADY           (),                              //                  .bready
		.f2h_ARID             (),                              //                  .arid
		.f2h_ARADDR           (),                              //                  .araddr
		.f2h_ARLEN            (),                              //                  .arlen
		.f2h_ARSIZE           (),                              //                  .arsize
		.f2h_ARBURST          (),                              //                  .arburst
		.f2h_ARLOCK           (),                              //                  .arlock
		.f2h_ARCACHE          (),                              //                  .arcache
		.f2h_ARPROT           (),                              //                  .arprot
		.f2h_ARVALID          (),                              //                  .arvalid
		.f2h_ARREADY          (),                              //                  .arready
		.f2h_ARUSER           (),                              //                  .aruser
		.f2h_RID              (),                              //                  .rid
		.f2h_RDATA            (),                              //                  .rdata
		.f2h_RRESP            (),                              //                  .rresp
		.f2h_RLAST            (),                              //                  .rlast
		.f2h_RVALID           (),                              //                  .rvalid
		.f2h_RREADY           (),                              //                  .rready
		.h2f_lw_axi_clk       (clk_clk),                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID          (hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR        (hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN         (hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE        (hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST       (hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK        (hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE       (hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT        (hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID       (hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY       (hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID           (hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA         (hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB         (hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST         (hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID        (hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY        (hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID           (hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP         (hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID        (hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY        (hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID          (hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR        (hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN         (hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE        (hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST       (hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK        (hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE       (hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT        (hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID       (hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY       (hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID           (hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA         (hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP         (hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST         (hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID        (hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY        (hps_h2f_lw_axi_master_rready)   //                  .rready
	);

	hps_gpio0 gpio0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_gpio0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio0_s1_readdata),   //                    .readdata
		.in_port    (gpio0_external_connection_in_port),     // external_connection.export
		.out_port   (gpio0_external_connection_out_port)     //                    .export
	);

	hps_gpio0 gpio1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_gpio1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio1_s1_readdata),   //                    .readdata
		.in_port    (gpio1_external_connection_in_port),     // external_connection.export
		.out_port   (gpio1_external_connection_out_port)     //                    .export
	);

	hps_keys keys (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_keys_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keys_s1_readdata), //                    .readdata
		.in_port  (keys_external_connection_export)     // external_connection.export
	);

	hps_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	hps_sw sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_external_connection_export)     // external_connection.export
	);

	hps_mm_interconnect_0 mm_interconnect_0 (
		.HPS_h2f_lw_axi_master_awid                                        (hps_h2f_lw_axi_master_awid),                 //                                       HPS_h2f_lw_axi_master.awid
		.HPS_h2f_lw_axi_master_awaddr                                      (hps_h2f_lw_axi_master_awaddr),               //                                                            .awaddr
		.HPS_h2f_lw_axi_master_awlen                                       (hps_h2f_lw_axi_master_awlen),                //                                                            .awlen
		.HPS_h2f_lw_axi_master_awsize                                      (hps_h2f_lw_axi_master_awsize),               //                                                            .awsize
		.HPS_h2f_lw_axi_master_awburst                                     (hps_h2f_lw_axi_master_awburst),              //                                                            .awburst
		.HPS_h2f_lw_axi_master_awlock                                      (hps_h2f_lw_axi_master_awlock),               //                                                            .awlock
		.HPS_h2f_lw_axi_master_awcache                                     (hps_h2f_lw_axi_master_awcache),              //                                                            .awcache
		.HPS_h2f_lw_axi_master_awprot                                      (hps_h2f_lw_axi_master_awprot),               //                                                            .awprot
		.HPS_h2f_lw_axi_master_awvalid                                     (hps_h2f_lw_axi_master_awvalid),              //                                                            .awvalid
		.HPS_h2f_lw_axi_master_awready                                     (hps_h2f_lw_axi_master_awready),              //                                                            .awready
		.HPS_h2f_lw_axi_master_wid                                         (hps_h2f_lw_axi_master_wid),                  //                                                            .wid
		.HPS_h2f_lw_axi_master_wdata                                       (hps_h2f_lw_axi_master_wdata),                //                                                            .wdata
		.HPS_h2f_lw_axi_master_wstrb                                       (hps_h2f_lw_axi_master_wstrb),                //                                                            .wstrb
		.HPS_h2f_lw_axi_master_wlast                                       (hps_h2f_lw_axi_master_wlast),                //                                                            .wlast
		.HPS_h2f_lw_axi_master_wvalid                                      (hps_h2f_lw_axi_master_wvalid),               //                                                            .wvalid
		.HPS_h2f_lw_axi_master_wready                                      (hps_h2f_lw_axi_master_wready),               //                                                            .wready
		.HPS_h2f_lw_axi_master_bid                                         (hps_h2f_lw_axi_master_bid),                  //                                                            .bid
		.HPS_h2f_lw_axi_master_bresp                                       (hps_h2f_lw_axi_master_bresp),                //                                                            .bresp
		.HPS_h2f_lw_axi_master_bvalid                                      (hps_h2f_lw_axi_master_bvalid),               //                                                            .bvalid
		.HPS_h2f_lw_axi_master_bready                                      (hps_h2f_lw_axi_master_bready),               //                                                            .bready
		.HPS_h2f_lw_axi_master_arid                                        (hps_h2f_lw_axi_master_arid),                 //                                                            .arid
		.HPS_h2f_lw_axi_master_araddr                                      (hps_h2f_lw_axi_master_araddr),               //                                                            .araddr
		.HPS_h2f_lw_axi_master_arlen                                       (hps_h2f_lw_axi_master_arlen),                //                                                            .arlen
		.HPS_h2f_lw_axi_master_arsize                                      (hps_h2f_lw_axi_master_arsize),               //                                                            .arsize
		.HPS_h2f_lw_axi_master_arburst                                     (hps_h2f_lw_axi_master_arburst),              //                                                            .arburst
		.HPS_h2f_lw_axi_master_arlock                                      (hps_h2f_lw_axi_master_arlock),               //                                                            .arlock
		.HPS_h2f_lw_axi_master_arcache                                     (hps_h2f_lw_axi_master_arcache),              //                                                            .arcache
		.HPS_h2f_lw_axi_master_arprot                                      (hps_h2f_lw_axi_master_arprot),               //                                                            .arprot
		.HPS_h2f_lw_axi_master_arvalid                                     (hps_h2f_lw_axi_master_arvalid),              //                                                            .arvalid
		.HPS_h2f_lw_axi_master_arready                                     (hps_h2f_lw_axi_master_arready),              //                                                            .arready
		.HPS_h2f_lw_axi_master_rid                                         (hps_h2f_lw_axi_master_rid),                  //                                                            .rid
		.HPS_h2f_lw_axi_master_rdata                                       (hps_h2f_lw_axi_master_rdata),                //                                                            .rdata
		.HPS_h2f_lw_axi_master_rresp                                       (hps_h2f_lw_axi_master_rresp),                //                                                            .rresp
		.HPS_h2f_lw_axi_master_rlast                                       (hps_h2f_lw_axi_master_rlast),                //                                                            .rlast
		.HPS_h2f_lw_axi_master_rvalid                                      (hps_h2f_lw_axi_master_rvalid),               //                                                            .rvalid
		.HPS_h2f_lw_axi_master_rready                                      (hps_h2f_lw_axi_master_rready),               //                                                            .rready
		.clk_0_clk_clk                                                     (clk_clk),                                    //                                                   clk_0_clk.clk
		.HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),         // HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.keys_reset_reset_bridge_in_reset_reset                            (rst_controller_reset_out_reset),             //                            keys_reset_reset_bridge_in_reset.reset
		.Arduino_io_s1_address                                             (mm_interconnect_0_arduino_io_s1_address),    //                                               Arduino_io_s1.address
		.Arduino_io_s1_write                                               (mm_interconnect_0_arduino_io_s1_write),      //                                                            .write
		.Arduino_io_s1_readdata                                            (mm_interconnect_0_arduino_io_s1_readdata),   //                                                            .readdata
		.Arduino_io_s1_writedata                                           (mm_interconnect_0_arduino_io_s1_writedata),  //                                                            .writedata
		.Arduino_io_s1_chipselect                                          (mm_interconnect_0_arduino_io_s1_chipselect), //                                                            .chipselect
		.gpio0_s1_address                                                  (mm_interconnect_0_gpio0_s1_address),         //                                                    gpio0_s1.address
		.gpio0_s1_write                                                    (mm_interconnect_0_gpio0_s1_write),           //                                                            .write
		.gpio0_s1_readdata                                                 (mm_interconnect_0_gpio0_s1_readdata),        //                                                            .readdata
		.gpio0_s1_writedata                                                (mm_interconnect_0_gpio0_s1_writedata),       //                                                            .writedata
		.gpio0_s1_chipselect                                               (mm_interconnect_0_gpio0_s1_chipselect),      //                                                            .chipselect
		.gpio1_s1_address                                                  (mm_interconnect_0_gpio1_s1_address),         //                                                    gpio1_s1.address
		.gpio1_s1_write                                                    (mm_interconnect_0_gpio1_s1_write),           //                                                            .write
		.gpio1_s1_readdata                                                 (mm_interconnect_0_gpio1_s1_readdata),        //                                                            .readdata
		.gpio1_s1_writedata                                                (mm_interconnect_0_gpio1_s1_writedata),       //                                                            .writedata
		.gpio1_s1_chipselect                                               (mm_interconnect_0_gpio1_s1_chipselect),      //                                                            .chipselect
		.keys_s1_address                                                   (mm_interconnect_0_keys_s1_address),          //                                                     keys_s1.address
		.keys_s1_readdata                                                  (mm_interconnect_0_keys_s1_readdata),         //                                                            .readdata
		.led_s1_address                                                    (mm_interconnect_0_led_s1_address),           //                                                      led_s1.address
		.led_s1_write                                                      (mm_interconnect_0_led_s1_write),             //                                                            .write
		.led_s1_readdata                                                   (mm_interconnect_0_led_s1_readdata),          //                                                            .readdata
		.led_s1_writedata                                                  (mm_interconnect_0_led_s1_writedata),         //                                                            .writedata
		.led_s1_chipselect                                                 (mm_interconnect_0_led_s1_chipselect),        //                                                            .chipselect
		.sw_s1_address                                                     (mm_interconnect_0_sw_s1_address),            //                                                       sw_s1.address
		.sw_s1_readdata                                                    (mm_interconnect_0_sw_s1_readdata)            //                                                            .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_h2f_reset_reset),           // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
